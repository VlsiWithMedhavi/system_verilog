module tb();

initial begin
	$display("\t#########");
	$display("\t#\t#");
	$display("\t#\t#");
	$display("\t#\t#");
	$display("\t#\t#");
	$display("\t#\t#");
	$display("#########################");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#\t\t\t#");
	$display("#########################");
end

endmodule
